module top(output [7:0] LED);
	assign LED[0] = 1'b1;
	assign LED[7:1] = 7'b0;
endmodule
